-- Dit is test 2