-- Dit is test 1